library verilog;
use verilog.vl_types.all;
entity lzw_FSK_vlg_tst is
end lzw_FSK_vlg_tst;
